module n_bit_multiplier #(parameter N = 4)
(
   ________ _______ [___:___] a, // Input 1
   ________ _______ [___:___] b, // Input 2
   ________ _______ [___:___] p  // Output Product: a*b
);
 
	// You got this! :)
 
endmodule
